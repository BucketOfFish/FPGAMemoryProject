localparam MEMNROWS = 16; // 16 words
localparam MEMNCOLS = 16; // each word is 16 bits long
localparam ROWINDEXBITS = 4;
localparam COLINDEXBITS = 4;
