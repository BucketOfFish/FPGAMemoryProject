localparam MEMORYDEPTH = 16; // 16 words
localparam WORDLENGTH = 16; // each word is 16 bits long
localparam WORDINDEXBITS = 4;
localparam LETTERINDEXBITS = 4;
localparam MAXBACKLOG = 100;