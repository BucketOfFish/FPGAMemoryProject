localparam MEMNROWS = 128;
localparam MEMNCOLS = 512;
localparam ROWINDEXBITS = 7;
localparam COLINDEXBITS = 9;
