localparam MEMNROWS_HNM = 128;
localparam MEMNCOLS_HNM = 512;
localparam MEMNROWS_HCM = 128*512;
localparam ROWINDEXBITS = 7;
localparam COLINDEXBITS = 9;
